module concat31(result, inp);
    input inp;
    output [31:0] result;
		
	or o1(result[0], inp, 0);
	or o2(result[1], 0, 0);
	or o3(result[2], 0, 0);
	or o4(result[3], 0, 0);
	or o5(result[4], 0, 0);
	or o6(result[5], 0, 0);
	or o7(result[6], 0, 0);
	or o8(result[7], 0, 0);
	or o9(result[8], 0, 0);
	or o10(result[9], 0, 0);
	or o11(result[10], 0, 0);
	or o12(result[11], 0, 0);
	or o13(result[12], 0, 0);
	or o14(result[13], 0, 0);
	or o15(result[14], 0, 0);
	or o16(result[15], 0, 0);
	or o17(result[16], 0, 0);
	or o18(result[17], 0, 0);
	or o19(result[18], 0, 0);
	or o20(result[19], 0, 0);
	or o21(result[20], 0, 0);
	or o22(result[21], 0, 0);
	or o23(result[22], 0, 0);
	or o24(result[23], 0, 0);
	or o25(result[24], 0, 0);
	or o26(result[25], 0, 0);
	or o27(result[26], 0, 0);
	or o28(result[27], 0, 0);
	or o29(result[28], 0, 0);
	or o30(result[29], 0, 0);
	or o31(result[30], 0, 0);
	or o32(result[31], 0, 0);

    
endmodule