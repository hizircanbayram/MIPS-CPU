module and_opr(res, a, b);
input [31:0] a, b;
output [31:0] res;

and AO0(res[0], a[0], b[0]),
	 AO1(res[1], a[1], b[1]),
	 AO2(res[2], a[2], b[2]),
	 AO3(res[3], a[3], b[3]),
	 AO4(res[4], a[4], b[4]),
	 AO5(res[5], a[5], b[5]),
	 AO6(res[6], a[6], b[6]),
	 AO7(res[7], a[7], b[7]),
	 AO8(res[8], a[8], b[8]),
	 AO9(res[9], a[9], b[9]),
	 AO10(res[10], a[10], b[10]),
	 AO11(res[11], a[11], b[11]),
	 AO12(res[12], a[12], b[12]),
	 AO13(res[13], a[13], b[13]),
	 AO14(res[14], a[14], b[14]),
	 AO15(res[15], a[15], b[15]),
	 AO16(res[16], a[16], b[16]),
	 AO17(res[17], a[17], b[17]),
	 AO18(res[18], a[18], b[18]),
	 AO19(res[19], a[19], b[19]),
	 AO20(res[20], a[20], b[20]),
	 AO21(res[21], a[21], b[21]),
	 AO22(res[22], a[22], b[22]),
	 AO23(res[23], a[23], b[23]),
	 AO24(res[24], a[24], b[24]),
	 AO25(res[25], a[25], b[25]),
	 AO26(res[26], a[26], b[26]),
	 AO27(res[27], a[27], b[27]),
	 AO28(res[28], a[28], b[28]),
	 AO29(res[29], a[29], b[29]),
	 AO30(res[30], a[30], b[30]),
	 AO31(res[31], a[31], b[31]);

endmodule